`timescale 1ns / 1ps

module testbench_500Hz;

    // Inputs
    reg clk, reset, clk_enable;
    reg signed [15:0] x;
    wire signed [15:0] y;
    // Instantiate the Unit Under Test (UUT)
    iir DUT(
     .clk(clk),
     .clk_enable(clk_enable),
     .reset(reset),
     .filter_in(x),
     .filter_out(y)
     );

    // Generate clock with 100ns period
    initial clk = 0;
    always #20833 clk = ~clk;


    // Initialize and pass sinusoidal input data of 2kHz with sampling frequency of 48kHz
    initial begin
        x = 16'b0;
        reset = 1;
        clk = 0;
        #100;
        reset = 0;
        #200;
        reset = 1;
        clk_enable = 1;
        #100;

        x = 0; #20833; // Sample(1)
    x = 699; #20833; // Sample(2)
    x = 1070; #20833; // Sample(3)
    x = 949; #20833; // Sample(4)
    x = 415; #20833; // Sample(5)
    x = -247; #20833; // Sample(6)
    x = -690; #20833; // Sample(7)
    x = -675; #20833; // Sample(8)
    x = -191; #20833; // Sample(9)
    x = 541; #20833; // Sample(10)
    x = 1176; #20833; // Sample(11)
    x = 1417; #20833; // Sample(12)
    x = 1161; #20833; // Sample(13)
    x = 554; #20833; // Sample(14)
    x = -86; #20833; // Sample(15)
    x = -425; #20833; // Sample(16)
    x = -278; #20833; // Sample(17)
    x = 298; #20833; // Sample(18)
    x = 1032; #20833; // Sample(19)
    x = 1576; #20833; // Sample(20)
    x = 1673; #20833; // Sample(21)
    x = 1290; #20833; // Sample(22)
    x = 630; #20833; // Sample(23)
    x = 33; #20833; // Sample(24)
    x = -191; #20833; // Sample(25)
    x = 80; #20833; // Sample(26)
    x = 722; #20833; // Sample(27)
    x = 1428; #20833; // Sample(28)
    x = 1857; #20833; // Sample(29)
    x = 1805; #20833; // Sample(30)
    x = 1307; #20833; // Sample(31)
    x = 617; #20833; // Sample(32)
    x = 85; #20833; // Sample(33)
    x = -18; #20833; // Sample(34)
    x = 364; #20833; // Sample(35)
    x = 1046; #20833; // Sample(36)
    x = 1695; #20833; // Sample(37)
    x = 1991; #20833; // Sample(38)
    x = 1790; #20833; // Sample(39)
    x = 1194; #20833; // Sample(40)
    x = 500; #20833; // Sample(41)
    x = 52; #20833; // Sample(42)
    x = 73; #20833; // Sample(43)
    x = 551; #20833; // Sample(44)
    x = 1247; #20833; // Sample(45)
    x = 1812; #20833; // Sample(46)
    x = 1964; #20833; // Sample(47)
    x = 1622; #20833; // Sample(48)
    x = 951; #20833; // Sample(49)
    x = 279; #20833; // Sample(50)
    x = -68; #20833; // Sample(51)
    x = 77; #20833; // Sample(52)
    x = 632; #20833; // Sample(53)
    x = 1315; #20833; // Sample(54)
    x = 1777; #20833; // Sample(55)
    x = 1778; #20833; // Sample(56)
    x = 1309; #20833; // Sample(57)
    x = 590; #20833; // Sample(58)
    x = -33; #20833; // Sample(59)
    x = -264; #20833; // Sample(60)
    x = 0; #20833; // Sample(61)
    x = 613; #20833; // Sample(62)
    x = 1258; #20833; // Sample(63)
    x = 1600; #20833; // Sample(64)
    x = 1454; #20833; // Sample(65)
    x = 877; #20833; // Sample(66)
    x = 140; #20833; // Sample(67)
    x = -408; #20833; // Sample(68)
    x = -512; #20833; // Sample(69)
    x = -137; #20833; // Sample(70)
    x = 513; #20833; // Sample(71)
    x = 1098; #20833; // Sample(72)
    x = 1309; #20833; // Sample(73)
    x = 1023; #20833; // Sample(74)
    x = 364; #20833; // Sample(75)
    x = -360; #20833; // Sample(76)
    x = -809; #20833; // Sample(77)
    x = -779; #20833; // Sample(78)
    x = -304; #20833; // Sample(79)
    x = 361; #20833; // Sample(80)
    x = 866; #20833; // Sample(81)
    x = 942; #20833; // Sample(82)
    x = 530; #20833; // Sample(83)
    x = -183; #20833; // Sample(84)
    x = -864; #20833; // Sample(85)
    x = -1193; #20833; // Sample(86)
    x = -1027; #20833; // Sample(87)
    x = -467; #20833; // Sample(88)
    x = 191; #20833; // Sample(89)
    x = 601; #20833; // Sample(90)
    x = 541; #20833; // Sample(91)
    x = 24; #20833; // Sample(92)
    x = -713; #20833; // Sample(93)
    x = -1320; #20833; // Sample(94)
    x = -1514; #20833; // Sample(95)
    x = -1215; #20833; // Sample(96)
    x = -588; #20833; // Sample(97)
    x = 40; #20833; // Sample(98)
    x = 342; #20833; // Sample(99)
    x = 153; #20833; // Sample(100)
    x = -448; #20833; // Sample(101)
    x = -1177; #20833; // Sample(102)
    x = -1684; #20833; // Sample(103)
    x = -1732; #20833; // Sample(104)
    x = -1309; #20833; // Sample(105)
    x = -636; #20833; // Sample(106)
    x = -59; #20833; // Sample(107)
    x = 125; #20833; // Sample(108)
    x = -184; #20833; // Sample(109)
    x = -843; #20833; // Sample(110)
    x = -1533; #20833; // Sample(111)
    x = -1919; #20833; // Sample(112)
    x = -1817; #20833; // Sample(113)
    x = -1284; #20833; // Sample(114)
    x = -590; #20833; // Sample(115)
    x = -84; #20833; // Sample(116)
    x = -22; #20833; // Sample(117)
    x = -437; #20833; // Sample(118)
    x = -1127; #20833; // Sample(119)
    x = -1751; #20833; // Sample(120)
    x = -2000; #20833; // Sample(121)
    x = -1751; #20833; // Sample(122)
    x = -1127; #20833; // Sample(123)
    x = -437; #20833; // Sample(124)
    x = -22; #20833; // Sample(125)
    x = -84; #20833; // Sample(126)
    x = -590; #20833; // Sample(127)
    x = -1284; #20833; // Sample(128)
    x = -1817; #20833; // Sample(129)
    x = -1919; #20833; // Sample(130)
    x = -1533; #20833; // Sample(131)
    x = -843; #20833; // Sample(132)
    x = -184; #20833; // Sample(133)
    x = 125; #20833; // Sample(134)
    x = -59; #20833; // Sample(135)
    x = -636; #20833; // Sample(136)
    x = -1309; #20833; // Sample(137)
    x = -1732; #20833; // Sample(138)
    x = -1684; #20833; // Sample(139)
    x = -1177; #20833; // Sample(140)
    x = -448; #20833; // Sample(141)
    x = 153; #20833; // Sample(142)
    x = 342; #20833; // Sample(143)
    x = 40; #20833; // Sample(144)
    x = -588; #20833; // Sample(145)
    x = -1215; #20833; // Sample(146)
    x = -1514; #20833; // Sample(147)
    x = -1320; #20833; // Sample(148)
    x = -713; #20833; // Sample(149)
    x = 24; #20833; // Sample(150)
    x = 541; #20833; // Sample(151)
    x = 601; #20833; // Sample(152)
    x = 191; #20833; // Sample(153)
    x = -467; #20833; // Sample(154)
    x = -1027; #20833; // Sample(155)
    x = -1193; #20833; // Sample(156)
    x = -864; #20833; // Sample(157)
    x = -183; #20833; // Sample(158)
    x = 530; #20833; // Sample(159)
    x = 942; #20833; // Sample(160)
    x = 866; #20833; // Sample(161)
    x = 361; #20833; // Sample(162)
    x = -304; #20833; // Sample(163)
    x = -779; #20833; // Sample(164)
    x = -809; #20833; // Sample(165)
    x = -360; #20833; // Sample(166)
    x = 364; #20833; // Sample(167)
    x = 1023; #20833; // Sample(168)
    x = 1309; #20833; // Sample(169)
    x = 1098; #20833; // Sample(170)
    x = 513; #20833; // Sample(171)
    x = -137; #20833; // Sample(172)
    x = -512; #20833; // Sample(173)
    x = -408; #20833; // Sample(174)
    x = 140; #20833; // Sample(175)
    x = 877; #20833; // Sample(176)
    x = 1454; #20833; // Sample(177)
    x = 1600; #20833; // Sample(178)
    x = 1258; #20833; // Sample(179)
    x = 613; #20833; // Sample(180)
    x = 0; #20833; // Sample(181)
    x = -264; #20833; // Sample(182)
    x = -33; #20833; // Sample(183)
    x = 590; #20833; // Sample(184)
    x = 1309; #20833; // Sample(185)
    x = 1778; #20833; // Sample(186)
    x = 1777; #20833; // Sample(187)
    x = 1315; #20833; // Sample(188)
    x = 632; #20833; // Sample(189)
    x = 77; #20833; // Sample(190)
    x = -68; #20833; // Sample(191)
    x = 279; #20833; // Sample(192)
    x = 951; #20833; // Sample(193)
    x = 1622; #20833; // Sample(194)
    x = 1964; #20833; // Sample(195)
    x = 1812; #20833; // Sample(196)
    x = 1247; #20833; // Sample(197)
    x = 551; #20833; // Sample(198)
    x = 73; #20833; // Sample(199)
    x = 52; #20833; // Sample(200)
    x = 500; #20833; // Sample(201)
    x = 1194; #20833; // Sample(202)
    x = 1790; #20833; // Sample(203)
    x = 1991; #20833; // Sample(204)
    x = 1695; #20833; // Sample(205)
    x = 1046; #20833; // Sample(206)
    x = 364; #20833; // Sample(207)
    x = -18; #20833; // Sample(208)
    x = 85; #20833; // Sample(209)
    x = 617; #20833; // Sample(210)
    x = 1307; #20833; // Sample(211)
    x = 1805; #20833; // Sample(212)
    x = 1857; #20833; // Sample(213)
    x = 1428; #20833; // Sample(214)
    x = 722; #20833; // Sample(215)
    x = 80; #20833; // Sample(216)
    x = -191; #20833; // Sample(217)
    x = 33; #20833; // Sample(218)
    x = 630; #20833; // Sample(219)
    x = 1290; #20833; // Sample(220)
    x = 1673; #20833; // Sample(221)
    x = 1576; #20833; // Sample(222)
    x = 1032; #20833; // Sample(223)
    x = 298; #20833; // Sample(224)
    x = -278; #20833; // Sample(225)
    x = -425; #20833; // Sample(226)
    x = -86; #20833; // Sample(227)
    x = 554; #20833; // Sample(228)
    x = 1161; #20833; // Sample(229)
    x = 1417; #20833; // Sample(230)
    x = 1176; #20833; // Sample(231)
    x = 541; #20833; // Sample(232)
    x = -191; #20833; // Sample(233)
    x = -675; #20833; // Sample(234)
    x = -690; #20833; // Sample(235)
    x = -247; #20833; // Sample(236)
    x = 415; #20833; // Sample(237)
    x = 949; #20833; // Sample(238)
    x = 1070; #20833; // Sample(239)
    x = 699; #20833; // Sample(240)
    x = 0; #20833; // Sample(241)
    x = -699; #20833; // Sample(242)
    x = -1070; #20833; // Sample(243)
    x = -949; #20833; // Sample(244)
    x = -415; #20833; // Sample(245)
    x = 247; #20833; // Sample(246)
    x = 690; #20833; // Sample(247)
    x = 675; #20833; // Sample(248)
    x = 191; #20833; // Sample(249)
    x = -541; #20833; // Sample(250)
    x = -1176; #20833; // Sample(251)
    x = -1417; #20833; // Sample(252)
    x = -1161; #20833; // Sample(253)
    x = -554; #20833; // Sample(254)
    x = 86; #20833; // Sample(255)
    x = 425; #20833; // Sample(256)
    x = 278; #20833; // Sample(257)
    x = -298; #20833; // Sample(258)
    x = -1032; #20833; // Sample(259)
    x = -1576; #20833; // Sample(260)
    x = -1673; #20833; // Sample(261)
    x = -1290; #20833; // Sample(262)
    x = -630; #20833; // Sample(263)
    x = -33; #20833; // Sample(264)
    x = 191; #20833; // Sample(265)
    x = -80; #20833; // Sample(266)
    x = -722; #20833; // Sample(267)
    x = -1428; #20833; // Sample(268)
    x = -1857; #20833; // Sample(269)
    x = -1805; #20833; // Sample(270)
    x = -1307; #20833; // Sample(271)
    x = -617; #20833; // Sample(272)
    x = -85; #20833; // Sample(273)
    x = 18; #20833; // Sample(274)
    x = -364; #20833; // Sample(275)
    x = -1046; #20833; // Sample(276)
    x = -1695; #20833; // Sample(277)
    x = -1991; #20833; // Sample(278)
    x = -1790; #20833; // Sample(279)
    x = -1194; #20833; // Sample(280)
    x = -500; #20833; // Sample(281)
    x = -52; #20833; // Sample(282)
    x = -73; #20833; // Sample(283)
    x = -551; #20833; // Sample(284)
    x = -1247; #20833; // Sample(285)
    x = -1812; #20833; // Sample(286)
    x = -1964; #20833; // Sample(287)
    x = -1622; #20833; // Sample(288)
    x = -951; #20833; // Sample(289)
    x = -279; #20833; // Sample(290)
    x = 68; #20833; // Sample(291)
    x = -77; #20833; // Sample(292)
    x = -632; #20833; // Sample(293)
    x = -1315; #20833; // Sample(294)
    x = -1777; #20833; // Sample(295)
    x = -1778; #20833; // Sample(296)
    x = -1309; #20833; // Sample(297)
    x = -590; #20833; // Sample(298)
    x = 33; #20833; // Sample(299)
    x = 264; #20833; // Sample(300)
    x = 0; #20833; // Sample(301)
    x = -613; #20833; // Sample(302)
    x = -1258; #20833; // Sample(303)
    x = -1600; #20833; // Sample(304)
    x = -1454; #20833; // Sample(305)
    x = -877; #20833; // Sample(306)
    x = -140; #20833; // Sample(307)
    x = 408; #20833; // Sample(308)
    x = 512; #20833; // Sample(309)
    x = 137; #20833; // Sample(310)
    x = -513; #20833; // Sample(311)
    x = -1098; #20833; // Sample(312)
    x = -1309; #20833; // Sample(313)
    x = -1023; #20833; // Sample(314)
    x = -364; #20833; // Sample(315)
    x = 360; #20833; // Sample(316)
    x = 809; #20833; // Sample(317)
    x = 779; #20833; // Sample(318)
    x = 304; #20833; // Sample(319)
    x = -361; #20833; // Sample(320)
    x = -866; #20833; // Sample(321)
    x = -942; #20833; // Sample(322)
    x = -530; #20833; // Sample(323)
    x = 183; #20833; // Sample(324)
    x = 864; #20833; // Sample(325)
    x = 1193; #20833; // Sample(326)
    x = 1027; #20833; // Sample(327)
    x = 467; #20833; // Sample(328)
    x = -191; #20833; // Sample(329)
    x = -601; #20833; // Sample(330)
    x = -541; #20833; // Sample(331)
    x = -24; #20833; // Sample(332)
    x = 713; #20833; // Sample(333)
    x = 1320; #20833; // Sample(334)
    x = 1514; #20833; // Sample(335)
    x = 1215; #20833; // Sample(336)
    x = 588; #20833; // Sample(337)
    x = -40; #20833; // Sample(338)
    x = -342; #20833; // Sample(339)
    x = -153; #20833; // Sample(340)
    x = 448; #20833; // Sample(341)
    x = 1177; #20833; // Sample(342)
    x = 1684; #20833; // Sample(343)
    x = 1732; #20833; // Sample(344)
    x = 1309; #20833; // Sample(345)
    x = 636; #20833; // Sample(346)
    x = 59; #20833; // Sample(347)
    x = -125; #20833; // Sample(348)
    x = 184; #20833; // Sample(349)
    x = 843; #20833; // Sample(350)
    x = 1533; #20833; // Sample(351)
    x = 1919; #20833; // Sample(352)
    x = 1817; #20833; // Sample(353)
    x = 1284; #20833; // Sample(354)
    x = 590; #20833; // Sample(355)
    x = 84; #20833; // Sample(356)
    x = 22; #20833; // Sample(357)
    x = 437; #20833; // Sample(358)
    x = 1127; #20833; // Sample(359)
    x = 1751; #20833; // Sample(360)
    x = 2000; #20833; // Sample(361)
    x = 1751; #20833; // Sample(362)
    x = 1127; #20833; // Sample(363)
    x = 437; #20833; // Sample(364)
    x = 22; #20833; // Sample(365)
    x = 84; #20833; // Sample(366)
    x = 590; #20833; // Sample(367)
    x = 1284; #20833; // Sample(368)
    x = 1817; #20833; // Sample(369)
    x = 1919; #20833; // Sample(370)
    x = 1533; #20833; // Sample(371)
    x = 843; #20833; // Sample(372)
    x = 184; #20833; // Sample(373)
    x = -125; #20833; // Sample(374)
    x = 59; #20833; // Sample(375)
    x = 636; #20833; // Sample(376)
    x = 1309; #20833; // Sample(377)
    x = 1732; #20833; // Sample(378)
    x = 1684; #20833; // Sample(379)
    x = 1177; #20833; // Sample(380)
    x = 448; #20833; // Sample(381)
    x = -153; #20833; // Sample(382)
    x = -342; #20833; // Sample(383)
    x = -40; #20833; // Sample(384)
    x = 588; #20833; // Sample(385)
    x = 1215; #20833; // Sample(386)
    x = 1514; #20833; // Sample(387)
    x = 1320; #20833; // Sample(388)
    x = 713; #20833; // Sample(389)
    x = -24; #20833; // Sample(390)
    x = -541; #20833; // Sample(391)
    x = -601; #20833; // Sample(392)
    x = -191; #20833; // Sample(393)
    x = 467; #20833; // Sample(394)
    x = 1027; #20833; // Sample(395)
    x = 1193; #20833; // Sample(396)
    x = 864; #20833; // Sample(397)
    x = 183; #20833; // Sample(398)
    x = -530; #20833; // Sample(399)
    x = -942; #20833; // Sample(400)
    x = -866; #20833; // Sample(401)
    x = -361; #20833; // Sample(402)
    x = 304; #20833; // Sample(403)
    x = 779; #20833; // Sample(404)
    x = 809; #20833; // Sample(405)
    x = 360; #20833; // Sample(406)
    x = -364; #20833; // Sample(407)
    x = -1023; #20833; // Sample(408)
    x = -1309; #20833; // Sample(409)
    x = -1098; #20833; // Sample(410)
    x = -513; #20833; // Sample(411)
    x = 137; #20833; // Sample(412)
    x = 512; #20833; // Sample(413)
    x = 408; #20833; // Sample(414)
    x = -140; #20833; // Sample(415)
    x = -877; #20833; // Sample(416)
    x = -1454; #20833; // Sample(417)
    x = -1600; #20833; // Sample(418)
    x = -1258; #20833; // Sample(419)
    x = -613; #20833; // Sample(420)
    x = 0; #20833; // Sample(421)
    x = 264; #20833; // Sample(422)
    x = 33; #20833; // Sample(423)
    x = -590; #20833; // Sample(424)
    x = -1309; #20833; // Sample(425)
    x = -1778; #20833; // Sample(426)
    x = -1777; #20833; // Sample(427)
    x = -1315; #20833; // Sample(428)
    x = -632; #20833; // Sample(429)
    x = -77; #20833; // Sample(430)
    x = 68; #20833; // Sample(431)
    x = -279; #20833; // Sample(432)
    x = -951; #20833; // Sample(433)
    x = -1622; #20833; // Sample(434)
    x = -1964; #20833; // Sample(435)
    x = -1812; #20833; // Sample(436)
    x = -1247; #20833; // Sample(437)
    x = -551; #20833; // Sample(438)
    x = -73; #20833; // Sample(439)
    x = -52; #20833; // Sample(440)
    x = -500; #20833; // Sample(441)
    x = -1194; #20833; // Sample(442)
    x = -1790; #20833; // Sample(443)
    x = -1991; #20833; // Sample(444)
    x = -1695; #20833; // Sample(445)
    x = -1046; #20833; // Sample(446)
    x = -364; #20833; // Sample(447)
    x = 18; #20833; // Sample(448)
    x = -85; #20833; // Sample(449)
    x = -617; #20833; // Sample(450)
    x = -1307; #20833; // Sample(451)
    x = -1805; #20833; // Sample(452)
    x = -1857; #20833; // Sample(453)
    x = -1428; #20833; // Sample(454)
    x = -722; #20833; // Sample(455)
    x = -80; #20833; // Sample(456)
    x = 191; #20833; // Sample(457)
    x = -33; #20833; // Sample(458)
    x = -630; #20833; // Sample(459)
    x = -1290; #20833; // Sample(460)
    x = -1673; #20833; // Sample(461)
    x = -1576; #20833; // Sample(462)
    x = -1032; #20833; // Sample(463)
    x = -298; #20833; // Sample(464)
    x = 278; #20833; // Sample(465)
    x = 425; #20833; // Sample(466)
    x = 86; #20833; // Sample(467)
    x = -554; #20833; // Sample(468)
    x = -1161; #20833; // Sample(469)
    x = -1417; #20833; // Sample(470)
    x = -1176; #20833; // Sample(471)
    x = -541; #20833; // Sample(472)
    x = 191; #20833; // Sample(473)
    x = 675; #20833; // Sample(474)
    x = 690; #20833; // Sample(475)
    x = 247; #20833; // Sample(476)
    x = -415; #20833; // Sample(477)
    x = -949; #20833; // Sample(478)
    x = -1070; #20833; // Sample(479)
    x = -699; #20833; // Sample(480)
    x = 0; #20833; // Sample(481)
    x = 699; #20833; // Sample(482)
    x = 1070; #20833; // Sample(483)
    x = 949; #20833; // Sample(484)
    x = 415; #20833; // Sample(485)
    x = -247; #20833; // Sample(486)
    x = -690; #20833; // Sample(487)
    x = -675; #20833; // Sample(488)
    x = -191; #20833; // Sample(489)
    x = 541; #20833; // Sample(490)
    x = 1176; #20833; // Sample(491)
    x = 1417; #20833; // Sample(492)
    x = 1161; #20833; // Sample(493)
    x = 554; #20833; // Sample(494)
    x = -86; #20833; // Sample(495)
    x = -425; #20833; // Sample(496)
    x = -278; #20833; // Sample(497)
    x = 298; #20833; // Sample(498)
    x = 1032; #20833; // Sample(499)
    x = 1576; #20833; // Sample(500)
    x = 1673; #20833; // Sample(501)
    x = 1290; #20833; // Sample(502)
    x = 630; #20833; // Sample(503)
    x = 33; #20833; // Sample(504)
    x = -191; #20833; // Sample(505)
    x = 80; #20833; // Sample(506)
    x = 722; #20833; // Sample(507)
    x = 1428; #20833; // Sample(508)
    x = 1857; #20833; // Sample(509)
    x = 1805; #20833; // Sample(510)
    x = 1307; #20833; // Sample(511)
    x = 617; #20833; // Sample(512)
    x = 85; #20833; // Sample(513)
    x = -18; #20833; // Sample(514)
    x = 364; #20833; // Sample(515)
    x = 1046; #20833; // Sample(516)
    x = 1695; #20833; // Sample(517)
    x = 1991; #20833; // Sample(518)
    x = 1790; #20833; // Sample(519)
    x = 1194; #20833; // Sample(520)
    x = 500; #20833; // Sample(521)
    x = 52; #20833; // Sample(522)
    x = 73; #20833; // Sample(523)
    x = 551; #20833; // Sample(524)
    x = 1247; #20833; // Sample(525)
    x = 1812; #20833; // Sample(526)
    x = 1964; #20833; // Sample(527)
    x = 1622; #20833; // Sample(528)
    x = 951; #20833; // Sample(529)
    x = 279; #20833; // Sample(530)
    x = -68; #20833; // Sample(531)
    x = 77; #20833; // Sample(532)
    x = 632; #20833; // Sample(533)
    x = 1315; #20833; // Sample(534)
    x = 1777; #20833; // Sample(535)
    x = 1778; #20833; // Sample(536)
    x = 1309; #20833; // Sample(537)
    x = 590; #20833; // Sample(538)
    x = -33; #20833; // Sample(539)
    x = -264; #20833; // Sample(540)
    x = 0; #20833; // Sample(541)
    x = 613; #20833; // Sample(542)
    x = 1258; #20833; // Sample(543)
    x = 1600; #20833; // Sample(544)
    x = 1454; #20833; // Sample(545)
    x = 877; #20833; // Sample(546)
    x = 140; #20833; // Sample(547)
    x = -408; #20833; // Sample(548)
    x = -512; #20833; // Sample(549)
    x = -137; #20833; // Sample(550)
    x = 513; #20833; // Sample(551)
    x = 1098; #20833; // Sample(552)
    x = 1309; #20833; // Sample(553)
    x = 1023; #20833; // Sample(554)
    x = 364; #20833; // Sample(555)
    x = -360; #20833; // Sample(556)
    x = -809; #20833; // Sample(557)
    x = -779; #20833; // Sample(558)
    x = -304; #20833; // Sample(559)
    x = 361; #20833; // Sample(560)
    x = 866; #20833; // Sample(561)
    x = 942; #20833; // Sample(562)
    x = 530; #20833; // Sample(563)
    x = -183; #20833; // Sample(564)
    x = -864; #20833; // Sample(565)
    x = -1193; #20833; // Sample(566)
    x = -1027; #20833; // Sample(567)
    x = -467; #20833; // Sample(568)
    x = 191; #20833; // Sample(569)
    x = 601; #20833; // Sample(570)
    x = 541; #20833; // Sample(571)
    x = 24; #20833; // Sample(572)
    x = -713; #20833; // Sample(573)
    x = -1320; #20833; // Sample(574)
    x = -1514; #20833; // Sample(575)
    x = -1215; #20833; // Sample(576)
    x = -588; #20833; // Sample(577)
    x = 40; #20833; // Sample(578)
    x = 342; #20833; // Sample(579)
    x = 153; #20833; // Sample(580)
    x = -448; #20833; // Sample(581)
    x = -1177; #20833; // Sample(582)
    x = -1684; #20833; // Sample(583)
    x = -1732; #20833; // Sample(584)
    x = -1309; #20833; // Sample(585)
    x = -636; #20833; // Sample(586)
    x = -59; #20833; // Sample(587)
    x = 125; #20833; // Sample(588)
    x = -184; #20833; // Sample(589)
    x = -843; #20833; // Sample(590)
    x = -1533; #20833; // Sample(591)
    x = -1919; #20833; // Sample(592)
    x = -1817; #20833; // Sample(593)
    x = -1284; #20833; // Sample(594)
    x = -590; #20833; // Sample(595)
    x = -84; #20833; // Sample(596)
    x = -22; #20833; // Sample(597)
    x = -437; #20833; // Sample(598)
    x = -1127; #20833; // Sample(599)
    x = -1751; #20833; // Sample(600)
    x = -2000; #20833; // Sample(601)
    x = -1751; #20833; // Sample(602)
    x = -1127; #20833; // Sample(603)
    x = -437; #20833; // Sample(604)
    x = -22; #20833; // Sample(605)
    x = -84; #20833; // Sample(606)
    x = -590; #20833; // Sample(607)
    x = -1284; #20833; // Sample(608)
    x = -1817; #20833; // Sample(609)
    x = -1919; #20833; // Sample(610)
    x = -1533; #20833; // Sample(611)
    x = -843; #20833; // Sample(612)
    x = -184; #20833; // Sample(613)
    x = 125; #20833; // Sample(614)
    x = -59; #20833; // Sample(615)
    x = -636; #20833; // Sample(616)
    x = -1309; #20833; // Sample(617)
    x = -1732; #20833; // Sample(618)
    x = -1684; #20833; // Sample(619)
    x = -1177; #20833; // Sample(620)
    x = -448; #20833; // Sample(621)
    x = 153; #20833; // Sample(622)
    x = 342; #20833; // Sample(623)
    x = 40; #20833; // Sample(624)
    x = -588; #20833; // Sample(625)
    x = -1215; #20833; // Sample(626)
    x = -1514; #20833; // Sample(627)
    x = -1320; #20833; // Sample(628)
    x = -713; #20833; // Sample(629)
    x = 24; #20833; // Sample(630)
    x = 541; #20833; // Sample(631)
    x = 601; #20833; // Sample(632)
    x = 191; #20833; // Sample(633)
    x = -467; #20833; // Sample(634)
    x = -1027; #20833; // Sample(635)
    x = -1193; #20833; // Sample(636)
    x = -864; #20833; // Sample(637)
    x = -183; #20833; // Sample(638)
    x = 530; #20833; // Sample(639)
    x = 942; #20833; // Sample(640)
    x = 866; #20833; // Sample(641)
    x = 361; #20833; // Sample(642)
    x = -304; #20833; // Sample(643)
    x = -779; #20833; // Sample(644)
    x = -809; #20833; // Sample(645)
    x = -360; #20833; // Sample(646)
    x = 364; #20833; // Sample(647)
    x = 1023; #20833; // Sample(648)
    x = 1309; #20833; // Sample(649)
    x = 1098; #20833; // Sample(650)
    x = 513; #20833; // Sample(651)
    x = -137; #20833; // Sample(652)
    x = -512; #20833; // Sample(653)
    x = -408; #20833; // Sample(654)
    x = 140; #20833; // Sample(655)
    x = 877; #20833; // Sample(656)
    x = 1454; #20833; // Sample(657)
    x = 1600; #20833; // Sample(658)
    x = 1258; #20833; // Sample(659)
    x = 613; #20833; // Sample(660)
    x = 0; #20833; // Sample(661)
    x = -264; #20833; // Sample(662)
    x = -33; #20833; // Sample(663)
    x = 590; #20833; // Sample(664)
    x = 1309; #20833; // Sample(665)
    x = 1778; #20833; // Sample(666)
    x = 1777; #20833; // Sample(667)
    x = 1315; #20833; // Sample(668)
    x = 632; #20833; // Sample(669)
    x = 77; #20833; // Sample(670)
    x = -68; #20833; // Sample(671)
    x = 279; #20833; // Sample(672)
    x = 951; #20833; // Sample(673)
    x = 1622; #20833; // Sample(674)
    x = 1964; #20833; // Sample(675)
    x = 1812; #20833; // Sample(676)
    x = 1247; #20833; // Sample(677)
    x = 551; #20833; // Sample(678)
    x = 73; #20833; // Sample(679)
    x = 52; #20833; // Sample(680)
    x = 500; #20833; // Sample(681)
    x = 1194; #20833; // Sample(682)
    x = 1790; #20833; // Sample(683)
    x = 1991; #20833; // Sample(684)
    x = 1695; #20833; // Sample(685)
    x = 1046; #20833; // Sample(686)
    x = 364; #20833; // Sample(687)
    x = -18; #20833; // Sample(688)
    x = 85; #20833; // Sample(689)
    x = 617; #20833; // Sample(690)
    x = 1307; #20833; // Sample(691)
    x = 1805; #20833; // Sample(692)
    x = 1857; #20833; // Sample(693)
    x = 1428; #20833; // Sample(694)
    x = 722; #20833; // Sample(695)
    x = 80; #20833; // Sample(696)
    x = -191; #20833; // Sample(697)
    x = 33; #20833; // Sample(698)
    x = 630; #20833; // Sample(699)
    x = 1290; #20833; // Sample(700)
    x = 1673; #20833; // Sample(701)
    x = 1576; #20833; // Sample(702)
    x = 1032; #20833; // Sample(703)
    x = 298; #20833; // Sample(704)
    x = -278; #20833; // Sample(705)
    x = -425; #20833; // Sample(706)
    x = -86; #20833; // Sample(707)
    x = 554; #20833; // Sample(708)
    x = 1161; #20833; // Sample(709)
    x = 1417; #20833; // Sample(710)
    x = 1176; #20833; // Sample(711)
    x = 541; #20833; // Sample(712)
    x = -191; #20833; // Sample(713)
    x = -675; #20833; // Sample(714)
    x = -690; #20833; // Sample(715)
    x = -247; #20833; // Sample(716)
    x = 415; #20833; // Sample(717)
    x = 949; #20833; // Sample(718)
    x = 1070; #20833; // Sample(719)
    x = 699; #20833; // Sample(720)
    x = 0; #20833; // Sample(721)
    x = -699; #20833; // Sample(722)
    x = -1070; #20833; // Sample(723)
    x = -949; #20833; // Sample(724)
    x = -415; #20833; // Sample(725)
    x = 247; #20833; // Sample(726)
    x = 690; #20833; // Sample(727)
    x = 675; #20833; // Sample(728)
    x = 191; #20833; // Sample(729)
    x = -541; #20833; // Sample(730)
    x = -1176; #20833; // Sample(731)
    x = -1417; #20833; // Sample(732)
    x = -1161; #20833; // Sample(733)
    x = -554; #20833; // Sample(734)
    x = 86; #20833; // Sample(735)
    x = 425; #20833; // Sample(736)
    x = 278; #20833; // Sample(737)
    x = -298; #20833; // Sample(738)
    x = -1032; #20833; // Sample(739)
    x = -1576; #20833; // Sample(740)
    x = -1673; #20833; // Sample(741)
    x = -1290; #20833; // Sample(742)
    x = -630; #20833; // Sample(743)
    x = -33; #20833; // Sample(744)
    x = 191; #20833; // Sample(745)
    x = -80; #20833; // Sample(746)
    x = -722; #20833; // Sample(747)
    x = -1428; #20833; // Sample(748)
    x = -1857; #20833; // Sample(749)
    x = -1805; #20833; // Sample(750)
    x = -1307; #20833; // Sample(751)
    x = -617; #20833; // Sample(752)
    x = -85; #20833; // Sample(753)
    x = 18; #20833; // Sample(754)
    x = -364; #20833; // Sample(755)
    x = -1046; #20833; // Sample(756)
    x = -1695; #20833; // Sample(757)
    x = -1991; #20833; // Sample(758)
    x = -1790; #20833; // Sample(759)
    x = -1194; #20833; // Sample(760)
    x = -500; #20833; // Sample(761)
    x = -52; #20833; // Sample(762)
    x = -73; #20833; // Sample(763)
    x = -551; #20833; // Sample(764)
    x = -1247; #20833; // Sample(765)
    x = -1812; #20833; // Sample(766)
    x = -1964; #20833; // Sample(767)
    x = -1622; #20833; // Sample(768)
    x = -951; #20833; // Sample(769)
    x = -279; #20833; // Sample(770)
    x = 68; #20833; // Sample(771)
    x = -77; #20833; // Sample(772)
    x = -632; #20833; // Sample(773)
    x = -1315; #20833; // Sample(774)
    x = -1777; #20833; // Sample(775)
    x = -1778; #20833; // Sample(776)
    x = -1309; #20833; // Sample(777)
    x = -590; #20833; // Sample(778)
    x = 33; #20833; // Sample(779)
    x = 264; #20833; // Sample(780)
    x = 0; #20833; // Sample(781)
    x = -613; #20833; // Sample(782)
    x = -1258; #20833; // Sample(783)
    x = -1600; #20833; // Sample(784)
    x = -1454; #20833; // Sample(785)
    x = -877; #20833; // Sample(786)
    x = -140; #20833; // Sample(787)
    x = 408; #20833; // Sample(788)
    x = 512; #20833; // Sample(789)
    x = 137; #20833; // Sample(790)
    x = -513; #20833; // Sample(791)
    x = -1098; #20833; // Sample(792)
    x = -1309; #20833; // Sample(793)
    x = -1023; #20833; // Sample(794)
    x = -364; #20833; // Sample(795)
    x = 360; #20833; // Sample(796)
    x = 809; #20833; // Sample(797)
    x = 779; #20833; // Sample(798)
    x = 304; #20833; // Sample(799)
    x = -361; #20833; // Sample(800)
    x = -866; #20833; // Sample(801)
    x = -942; #20833; // Sample(802)
    x = -530; #20833; // Sample(803)
    x = 183; #20833; // Sample(804)
    x = 864; #20833; // Sample(805)
    x = 1193; #20833; // Sample(806)
    x = 1027; #20833; // Sample(807)
    x = 467; #20833; // Sample(808)
    x = -191; #20833; // Sample(809)
    x = -601; #20833; // Sample(810)
    x = -541; #20833; // Sample(811)
    x = -24; #20833; // Sample(812)
    x = 713; #20833; // Sample(813)
    x = 1320; #20833; // Sample(814)
    x = 1514; #20833; // Sample(815)
    x = 1215; #20833; // Sample(816)
    x = 588; #20833; // Sample(817)
    x = -40; #20833; // Sample(818)
    x = -342; #20833; // Sample(819)
    x = -153; #20833; // Sample(820)
    x = 448; #20833; // Sample(821)
    x = 1177; #20833; // Sample(822)
    x = 1684; #20833; // Sample(823)
    x = 1732; #20833; // Sample(824)
    x = 1309; #20833; // Sample(825)
    x = 636; #20833; // Sample(826)
    x = 59; #20833; // Sample(827)
    x = -125; #20833; // Sample(828)
    x = 184; #20833; // Sample(829)
    x = 843; #20833; // Sample(830)
    x = 1533; #20833; // Sample(831)
    x = 1919; #20833; // Sample(832)
    x = 1817; #20833; // Sample(833)
    x = 1284; #20833; // Sample(834)
    x = 590; #20833; // Sample(835)
    x = 84; #20833; // Sample(836)
    x = 22; #20833; // Sample(837)
    x = 437; #20833; // Sample(838)
    x = 1127; #20833; // Sample(839)
    x = 1751; #20833; // Sample(840)
    x = 2000; #20833; // Sample(841)
    x = 1751; #20833; // Sample(842)
    x = 1127; #20833; // Sample(843)
    x = 437; #20833; // Sample(844)
    x = 22; #20833; // Sample(845)
    x = 84; #20833; // Sample(846)
    x = 590; #20833; // Sample(847)
    x = 1284; #20833; // Sample(848)
    x = 1817; #20833; // Sample(849)
    x = 1919; #20833; // Sample(850)
    x = 1533; #20833; // Sample(851)
    x = 843; #20833; // Sample(852)
    x = 184; #20833; // Sample(853)
    x = -125; #20833; // Sample(854)
    x = 59; #20833; // Sample(855)
    x = 636; #20833; // Sample(856)
    x = 1309; #20833; // Sample(857)
    x = 1732; #20833; // Sample(858)
    x = 1684; #20833; // Sample(859)
    x = 1177; #20833; // Sample(860)
    x = 448; #20833; // Sample(861)
    x = -153; #20833; // Sample(862)
    x = -342; #20833; // Sample(863)
    x = -40; #20833; // Sample(864)
    x = 588; #20833; // Sample(865)
    x = 1215; #20833; // Sample(866)
    x = 1514; #20833; // Sample(867)
    x = 1320; #20833; // Sample(868)
    x = 713; #20833; // Sample(869)
    x = -24; #20833; // Sample(870)
    x = -541; #20833; // Sample(871)
    x = -601; #20833; // Sample(872)
    x = -191; #20833; // Sample(873)
    x = 467; #20833; // Sample(874)
    x = 1027; #20833; // Sample(875)
    x = 1193; #20833; // Sample(876)
    x = 864; #20833; // Sample(877)
    x = 183; #20833; // Sample(878)
    x = -530; #20833; // Sample(879)
    x = -942; #20833; // Sample(880)
    x = -866; #20833; // Sample(881)
    x = -361; #20833; // Sample(882)
    x = 304; #20833; // Sample(883)
    x = 779; #20833; // Sample(884)
    x = 809; #20833; // Sample(885)
    x = 360; #20833; // Sample(886)
    x = -364; #20833; // Sample(887)
    x = -1023; #20833; // Sample(888)
    x = -1309; #20833; // Sample(889)
    x = -1098; #20833; // Sample(890)
    x = -513; #20833; // Sample(891)
    x = 137; #20833; // Sample(892)
    x = 512; #20833; // Sample(893)
    x = 408; #20833; // Sample(894)
    x = -140; #20833; // Sample(895)
    x = -877; #20833; // Sample(896)
    x = -1454; #20833; // Sample(897)
    x = -1600; #20833; // Sample(898)
    x = -1258; #20833; // Sample(899)
    x = -613; #20833; // Sample(900)
    x = 0; #20833; // Sample(901)
    x = 264; #20833; // Sample(902)
    x = 33; #20833; // Sample(903)
    x = -590; #20833; // Sample(904)
    x = -1309; #20833; // Sample(905)
    x = -1778; #20833; // Sample(906)
    x = -1777; #20833; // Sample(907)
    x = -1315; #20833; // Sample(908)
    x = -632; #20833; // Sample(909)
    x = -77; #20833; // Sample(910)
    x = 68; #20833; // Sample(911)
    x = -279; #20833; // Sample(912)
    x = -951; #20833; // Sample(913)
    x = -1622; #20833; // Sample(914)
    x = -1964; #20833; // Sample(915)
    x = -1812; #20833; // Sample(916)
    x = -1247; #20833; // Sample(917)
    x = -551; #20833; // Sample(918)
    x = -73; #20833; // Sample(919)
    x = -52; #20833; // Sample(920)
    x = -500; #20833; // Sample(921)
    x = -1194; #20833; // Sample(922)
    x = -1790; #20833; // Sample(923)
    x = -1991; #20833; // Sample(924)
    x = -1695; #20833; // Sample(925)
    x = -1046; #20833; // Sample(926)
    x = -364; #20833; // Sample(927)
    x = 18; #20833; // Sample(928)
    x = -85; #20833; // Sample(929)
    x = -617; #20833; // Sample(930)
    x = -1307; #20833; // Sample(931)
    x = -1805; #20833; // Sample(932)
    x = -1857; #20833; // Sample(933)
    x = -1428; #20833; // Sample(934)
    x = -722; #20833; // Sample(935)
    x = -80; #20833; // Sample(936)
    x = 191; #20833; // Sample(937)
    x = -33; #20833; // Sample(938)
    x = -630; #20833; // Sample(939)
    x = -1290; #20833; // Sample(940)
    x = -1673; #20833; // Sample(941)
    x = -1576; #20833; // Sample(942)
    x = -1032; #20833; // Sample(943)
    x = -298; #20833; // Sample(944)
    x = 278; #20833; // Sample(945)
    x = 425; #20833; // Sample(946)
    x = 86; #20833; // Sample(947)
    x = -554; #20833; // Sample(948)
    x = -1161; #20833; // Sample(949)
    x = -1417; #20833; // Sample(950)
    x = -1176; #20833; // Sample(951)
    x = -541; #20833; // Sample(952)
    x = 191; #20833; // Sample(953)
    x = 675; #20833; // Sample(954)
    x = 690; #20833; // Sample(955)
    x = 247; #20833; // Sample(956)
    x = -415; #20833; // Sample(957)
    x = -949; #20833; // Sample(958)
    x = -1070; #20833; // Sample(959)
    x = -699; #20833; // Sample(960)
    x = 0; #20833; // Sample(961)
    x = 699; #20833; // Sample(962)
    x = 1070; #20833; // Sample(963)
    x = 949; #20833; // Sample(964)
    x = 415; #20833; // Sample(965)
    x = -247; #20833; // Sample(966)
    x = -690; #20833; // Sample(967)
    x = -675; #20833; // Sample(968)
    x = -191; #20833; // Sample(969)
    x = 541; #20833; // Sample(970)
    x = 1176; #20833; // Sample(971)
    x = 1417; #20833; // Sample(972)
    x = 1161; #20833; // Sample(973)
    x = 554; #20833; // Sample(974)
    x = -86; #20833; // Sample(975)
    x = -425; #20833; // Sample(976)
    x = -278; #20833; // Sample(977)
    x = 298; #20833; // Sample(978)
    x = 1032; #20833; // Sample(979)
    x = 1576; #20833; // Sample(980)
    x = 1673; #20833; // Sample(981)
    x = 1290; #20833; // Sample(982)
    x = 630; #20833; // Sample(983)
    x = 33; #20833; // Sample(984)
    x = -191; #20833; // Sample(985)
    x = 80; #20833; // Sample(986)
    x = 722; #20833; // Sample(987)
    x = 1428; #20833; // Sample(988)
    x = 1857; #20833; // Sample(989)
    x = 1805; #20833; // Sample(990)
    x = 1307; #20833; // Sample(991)
    x = 617; #20833; // Sample(992)
    x = 85; #20833; // Sample(993)
    x = -18; #20833; // Sample(994)
    x = 364; #20833; // Sample(995)
    x = 1046; #20833; // Sample(996)
    x = 1695; #20833; // Sample(997)
    x = 1991; #20833; // Sample(998)
    x = 1790; #20833; // Sample(999)
    x = 1194; #20833; // Sample(1000)
        $stop;
    end
endmodule
