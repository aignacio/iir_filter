`timescale 1ns / 1ps

module testbench_500Hz;

    // Inputs
    reg clk, reset;
    reg signed [31:0] x;
    wire signed [31:0] y;
    // Instantiate the Unit Under Test (UUT)
    iir DUT(
      .clk(clk),
      .rst(reset),
      .x(x),
      .y(y)
    );

    // Generate clock with 100ns period
    initial clk = 0;
    always #20833 clk = ~clk;

    initial begin
        x = 32'd0;
        reset = 1;
        clk = 0;
        #10;
        reset = 0;
        #20;
        reset = 1;
        #10;
        x =               67; #20833; // Sample(1)
        x =             -456; #20833; // Sample(2)
        x =               19; #20833; // Sample(3)
        x =               28; #20833; // Sample(4)
        x =              160; #20833; // Sample(5)
        x =               39; #20833; // Sample(6)
        x =              142; #20833; // Sample(7)
        x =              151; #20833; // Sample(8)
        x =              117; #20833; // Sample(9)
        x =              294; #20833; // Sample(10)
        x =              199; #20833; // Sample(11)
        x =              363; #20833; // Sample(12)
        x =              100; #20833; // Sample(13)
        x =              525; #20833; // Sample(14)
        x =               78; #20833; // Sample(15)
        x =              195; #20833; // Sample(16)
        x =              -19; #20833; // Sample(17)
        x =              147; #20833; // Sample(18)
        x =              515; #20833; // Sample(19)
        x =              373; #20833; // Sample(20)
        x =              110; #20833; // Sample(21)
        x =              389; #20833; // Sample(22)
        x =              161; #20833; // Sample(23)
        x =              -98; #20833; // Sample(24)
        x =              198; #20833; // Sample(25)
        x =              673; #20833; // Sample(26)
        x =              338; #20833; // Sample(27)
        x =              -79; #20833; // Sample(28)
        x =              424; #20833; // Sample(29)
        x =              653; #20833; // Sample(30)
        x =              269; #20833; // Sample(31)
        x =              241; #20833; // Sample(32)
        x =              374; #20833; // Sample(33)
        x =               92; #20833; // Sample(34)
        x =              296; #20833; // Sample(35)
        x =              707; #20833; // Sample(36)
        x =               46; #20833; // Sample(37)
        x =              212; #20833; // Sample(38)
        x =              262; #20833; // Sample(39)
        x =              251; #20833; // Sample(40)
        x =              315; #20833; // Sample(41)
        x =               94; #20833; // Sample(42)
        x =              -26; #20833; // Sample(43)
        x =               84; #20833; // Sample(44)
        x =             -286; #20833; // Sample(45)
        x =               18; #20833; // Sample(46)
        x =              459; #20833; // Sample(47)
        x =              -86; #20833; // Sample(48)
        x =               70; #20833; // Sample(49)
        x =               77; #20833; // Sample(50)
        x =               38; #20833; // Sample(51)
        x =              -44; #20833; // Sample(52)
        x =             -200; #20833; // Sample(53)
        x =              -27; #20833; // Sample(54)
        x =              -67; #20833; // Sample(55)
        x =             -100; #20833; // Sample(56)
        x =              -33; #20833; // Sample(57)
        x =             -199; #20833; // Sample(58)
        x =             -407; #20833; // Sample(59)
        x =             -343; #20833; // Sample(60)
        x =              -78; #20833; // Sample(61)
        x =              -28; #20833; // Sample(62)
        x =             -358; #20833; // Sample(63)
        x =             -503; #20833; // Sample(64)
        x =             -454; #20833; // Sample(65)
        x =              -75; #20833; // Sample(66)
        x =             -101; #20833; // Sample(67)
        x =             -133; #20833; // Sample(68)
        x =             -103; #20833; // Sample(69)
        x =             -299; #20833; // Sample(70)
        x =             -267; #20833; // Sample(71)
        x =             -161; #20833; // Sample(72)
        x =             -123; #20833; // Sample(73)
        x =              191; #20833; // Sample(74)
        x =             -482; #20833; // Sample(75)
        x =             -272; #20833; // Sample(76)
        x =             -206; #20833; // Sample(77)
        x =             -506; #20833; // Sample(78)
        x =             -562; #20833; // Sample(79)
        x =             -238; #20833; // Sample(80)
        x =             -396; #20833; // Sample(81)
        x =             -249; #20833; // Sample(82)
        x =             -421; #20833; // Sample(83)
        x =             -245; #20833; // Sample(84)
        x =             -193; #20833; // Sample(85)
        x =             -624; #20833; // Sample(86)
        x =              -37; #20833; // Sample(87)
        x =             -554; #20833; // Sample(88)
        x =             -101; #20833; // Sample(89)
        x =             -129; #20833; // Sample(90)
        x =              -70; #20833; // Sample(91)
        x =              197; #20833; // Sample(92)
        x =             -374; #20833; // Sample(93)
        x =             -191; #20833; // Sample(94)
        x =             -186; #20833; // Sample(95)
        x =              278; #20833; // Sample(96)
        x =              253; #20833; // Sample(97)
        x =              156; #20833; // Sample(98)
        x =             -260; #20833; // Sample(99)
        x =              -30; #20833; // Sample(100)
        x =              179; #20833; // Sample(101)
        x =              164; #20833; // Sample(102)
        x =              -10; #20833; // Sample(103)
        x =              423; #20833; // Sample(104)
        x =               39; #20833; // Sample(105)
        x =              241; #20833; // Sample(106)
        x =              568; #20833; // Sample(107)
        x =              532; #20833; // Sample(108)
        x =              174; #20833; // Sample(109)
        x =              371; #20833; // Sample(110)
        x =              562; #20833; // Sample(111)
        x =               66; #20833; // Sample(112)
        x =              445; #20833; // Sample(113)
        x =              628; #20833; // Sample(114)
        x =              471; #20833; // Sample(115)
        x =              522; #20833; // Sample(116)
        x =              290; #20833; // Sample(117)
        x =               47; #20833; // Sample(118)
        x =              157; #20833; // Sample(119)
        x =              597; #20833; // Sample(120)
        x =              314; #20833; // Sample(121)
        x =              458; #20833; // Sample(122)
        x =              102; #20833; // Sample(123)
        x =              -47; #20833; // Sample(124)
        x =             -105; #20833; // Sample(125)
        x =              338; #20833; // Sample(126)
        x =             -133; #20833; // Sample(127)
        x =              543; #20833; // Sample(128)
        x =              479; #20833; // Sample(129)
        x =              307; #20833; // Sample(130)
        x =              435; #20833; // Sample(131)
        x =              206; #20833; // Sample(132)
        x =             -133; #20833; // Sample(133)
        x =              174; #20833; // Sample(134)
        x =               55; #20833; // Sample(135)
        x =              405; #20833; // Sample(136)
        x =              216; #20833; // Sample(137)
        x =              211; #20833; // Sample(138)
        x =               45; #20833; // Sample(139)
        x =              -72; #20833; // Sample(140)
        x =              131; #20833; // Sample(141)
        x =              -23; #20833; // Sample(142)
        x =              301; #20833; // Sample(143)
        x =              -49; #20833; // Sample(144)
        x =             -150; #20833; // Sample(145)
        x =              -61; #20833; // Sample(146)
        x =              165; #20833; // Sample(147)
        x =             -166; #20833; // Sample(148)
        x =              -96; #20833; // Sample(149)
        x =             -374; #20833; // Sample(150)
        x =              -92; #20833; // Sample(151)
        x =             -205; #20833; // Sample(152)
        x =             -234; #20833; // Sample(153)
        x =             -140; #20833; // Sample(154)
        x =             -178; #20833; // Sample(155)
        x =             -198; #20833; // Sample(156)
        x =              354; #20833; // Sample(157)
        x =              -29; #20833; // Sample(158)
        x =               80; #20833; // Sample(159)
        x =               65; #20833; // Sample(160)
        x =             -314; #20833; // Sample(161)
        x =             -361; #20833; // Sample(162)
        x =             -591; #20833; // Sample(163)
        x =             -467; #20833; // Sample(164)
        x =             -344; #20833; // Sample(165)
        x =             -311; #20833; // Sample(166)
        x =             -236; #20833; // Sample(167)
        x =             -270; #20833; // Sample(168)
        x =             -525; #20833; // Sample(169)
        x =             -361; #20833; // Sample(170)
        x =               30; #20833; // Sample(171)
        x =             -351; #20833; // Sample(172)
        x =             -464; #20833; // Sample(173)
        x =             -332; #20833; // Sample(174)
        x =             -214; #20833; // Sample(175)
        x =             -342; #20833; // Sample(176)
        x =             -341; #20833; // Sample(177)
        x =             -314; #20833; // Sample(178)
        x =              -13; #20833; // Sample(179)
        x =              -67; #20833; // Sample(180)
        x =             -354; #20833; // Sample(181)
        x =             -339; #20833; // Sample(182)
        x =             -512; #20833; // Sample(183)
        x =               46; #20833; // Sample(184)
        x =             -170; #20833; // Sample(185)
        x =             -179; #20833; // Sample(186)
        x =              -81; #20833; // Sample(187)
        x =             -342; #20833; // Sample(188)
        x =             -252; #20833; // Sample(189)
        x =              -24; #20833; // Sample(190)
        x =             -100; #20833; // Sample(191)
        x =             -409; #20833; // Sample(192)
        x =             -146; #20833; // Sample(193)
        x =               70; #20833; // Sample(194)
        x =              242; #20833; // Sample(195)
        x =               76; #20833; // Sample(196)
        x =              105; #20833; // Sample(197)
        x =                5; #20833; // Sample(198)
        x =              155; #20833; // Sample(199)
        x =              236; #20833; // Sample(200)
        x =              -21; #20833; // Sample(201)
        x =              366; #20833; // Sample(202)
        x =             -132; #20833; // Sample(203)
        x =              189; #20833; // Sample(204)
        x =              168; #20833; // Sample(205)
        x =              538; #20833; // Sample(206)
        x =              179; #20833; // Sample(207)
        x =              861; #20833; // Sample(208)
        x =              208; #20833; // Sample(209)
        x =              133; #20833; // Sample(210)
        x =              718; #20833; // Sample(211)
        x =              280; #20833; // Sample(212)
        x =              241; #20833; // Sample(213)
        x =              322; #20833; // Sample(214)
        x =              107; #20833; // Sample(215)
        x =               22; #20833; // Sample(216)
        x =              178; #20833; // Sample(217)
        x =              312; #20833; // Sample(218)
        x =              514; #20833; // Sample(219)
        x =              524; #20833; // Sample(220)
        x =              381; #20833; // Sample(221)
        x =              511; #20833; // Sample(222)
        x =              775; #20833; // Sample(223)
        x =              393; #20833; // Sample(224)
        x =              443; #20833; // Sample(225)
        x =              192; #20833; // Sample(226)
        x =              466; #20833; // Sample(227)
        x =               12; #20833; // Sample(228)
        x =              149; #20833; // Sample(229)
        x =               35; #20833; // Sample(230)
        x =               77; #20833; // Sample(231)
        x =              545; #20833; // Sample(232)
        x =              111; #20833; // Sample(233)
        x =               52; #20833; // Sample(234)
        x =              311; #20833; // Sample(235)
        x =               36; #20833; // Sample(236)
        x =              139; #20833; // Sample(237)
        x =              164; #20833; // Sample(238)
        x =             -126; #20833; // Sample(239)
        x =              -47; #20833; // Sample(240)
        x =              365; #20833; // Sample(241)
        x =                6; #20833; // Sample(242)
        x =              133; #20833; // Sample(243)
        x =              184; #20833; // Sample(244)
        x =               32; #20833; // Sample(245)
        x =              -72; #20833; // Sample(246)
        x =              129; #20833; // Sample(247)
        x =             -372; #20833; // Sample(248)
        x =               80; #20833; // Sample(249)
        x =             -567; #20833; // Sample(250)
        x =             -423; #20833; // Sample(251)
        x =             -279; #20833; // Sample(252)
        x =             -228; #20833; // Sample(253)
        x =             -536; #20833; // Sample(254)
        x =              -90; #20833; // Sample(255)
        x =             -264; #20833; // Sample(256)
        x =             -469; #20833; // Sample(257)
        x =             -496; #20833; // Sample(258)
        x =             -460; #20833; // Sample(259)
        x =             -443; #20833; // Sample(260)
        x =             -314; #20833; // Sample(261)
        x =             -304; #20833; // Sample(262)
        x =             -408; #20833; // Sample(263)
        x =             -315; #20833; // Sample(264)
        x =             -423; #20833; // Sample(265)
        x =             -265; #20833; // Sample(266)
        x =               -2; #20833; // Sample(267)
        x =             -130; #20833; // Sample(268)
        x =             -368; #20833; // Sample(269)
        x =             -256; #20833; // Sample(270)
        x =             -307; #20833; // Sample(271)
        x =             -350; #20833; // Sample(272)
        x =             -320; #20833; // Sample(273)
        x =              -38; #20833; // Sample(274)
        x =             -342; #20833; // Sample(275)
        x =             -190; #20833; // Sample(276)
        x =              -95; #20833; // Sample(277)
        x =             -395; #20833; // Sample(278)
        x =             -470; #20833; // Sample(279)
        x =              -21; #20833; // Sample(280)
        x =              -77; #20833; // Sample(281)
        x =             -235; #20833; // Sample(282)
        x =              100; #20833; // Sample(283)
        x =              -36; #20833; // Sample(284)
        x =             -155; #20833; // Sample(285)
        x =             -143; #20833; // Sample(286)
        x =             -134; #20833; // Sample(287)
        x =             -228; #20833; // Sample(288)
        x =              519; #20833; // Sample(289)
        x =             -412; #20833; // Sample(290)
        x =               91; #20833; // Sample(291)
        x =               60; #20833; // Sample(292)
        x =             -166; #20833; // Sample(293)
        x =               68; #20833; // Sample(294)
        x =              189; #20833; // Sample(295)
        x =              328; #20833; // Sample(296)
        x =              171; #20833; // Sample(297)
        x =              278; #20833; // Sample(298)
        x =              516; #20833; // Sample(299)
        x =              177; #20833; // Sample(300)
        x =              103; #20833; // Sample(301)
        x =              -46; #20833; // Sample(302)
        x =              399; #20833; // Sample(303)
        x =              152; #20833; // Sample(304)
        x =              530; #20833; // Sample(305)
        x =              283; #20833; // Sample(306)
        x =              251; #20833; // Sample(307)
        x =              177; #20833; // Sample(308)
        x =              192; #20833; // Sample(309)
        x =               54; #20833; // Sample(310)
        x =              411; #20833; // Sample(311)
        x =              219; #20833; // Sample(312)
        x =              421; #20833; // Sample(313)
        x =              -22; #20833; // Sample(314)
        x =              362; #20833; // Sample(315)
        x =              120; #20833; // Sample(316)
        x =               -7; #20833; // Sample(317)
        x =              239; #20833; // Sample(318)
        x =              394; #20833; // Sample(319)
        x =              465; #20833; // Sample(320)
        x =              494; #20833; // Sample(321)
        x =              177; #20833; // Sample(322)
        x =               56; #20833; // Sample(323)
        x =              802; #20833; // Sample(324)
        x =              108; #20833; // Sample(325)
        x =               64; #20833; // Sample(326)
        x =              273; #20833; // Sample(327)
        x =              -37; #20833; // Sample(328)
        x =               24; #20833; // Sample(329)
        x =             -156; #20833; // Sample(330)
        x =               77; #20833; // Sample(331)
        x =             -117; #20833; // Sample(332)
        x =              152; #20833; // Sample(333)
        x =               95; #20833; // Sample(334)
        x =              -97; #20833; // Sample(335)
        x =              -53; #20833; // Sample(336)
        x =             -108; #20833; // Sample(337)
        x =               12; #20833; // Sample(338)
        x =             -163; #20833; // Sample(339)
        x =               -8; #20833; // Sample(340)
        x =             -239; #20833; // Sample(341)
        x =               15; #20833; // Sample(342)
        x =             -146; #20833; // Sample(343)
        x =             -521; #20833; // Sample(344)
        x =             -114; #20833; // Sample(345)
        x =               12; #20833; // Sample(346)
        x =               56; #20833; // Sample(347)
        x =             -155; #20833; // Sample(348)
        x =               68; #20833; // Sample(349)
        x =              -95; #20833; // Sample(350)
        x =              160; #20833; // Sample(351)
        x =             -199; #20833; // Sample(352)
        x =             -169; #20833; // Sample(353)
        x =             -187; #20833; // Sample(354)
        x =             -172; #20833; // Sample(355)
        x =             -127; #20833; // Sample(356)
        x =              -89; #20833; // Sample(357)
        x =             -480; #20833; // Sample(358)
        x =             -542; #20833; // Sample(359)
        x =              -47; #20833; // Sample(360)
        x =             -117; #20833; // Sample(361)
        x =             -459; #20833; // Sample(362)
        x =             -306; #20833; // Sample(363)
        x =               55; #20833; // Sample(364)
        x =             -508; #20833; // Sample(365)
        x =             -222; #20833; // Sample(366)
        x =             -539; #20833; // Sample(367)
        x =             -236; #20833; // Sample(368)
        x =             -202; #20833; // Sample(369)
        x =             -283; #20833; // Sample(370)
        x =              -60; #20833; // Sample(371)
        x =             -252; #20833; // Sample(372)
        x =               12; #20833; // Sample(373)
        x =                9; #20833; // Sample(374)
        x =             -235; #20833; // Sample(375)
        x =             -118; #20833; // Sample(376)
        x =             -110; #20833; // Sample(377)
        x =               50; #20833; // Sample(378)
        x =              120; #20833; // Sample(379)
        x =               54; #20833; // Sample(380)
        x =              -73; #20833; // Sample(381)
        x =             -227; #20833; // Sample(382)
        x =             -282; #20833; // Sample(383)
        x =              188; #20833; // Sample(384)
        x =              377; #20833; // Sample(385)
        x =               71; #20833; // Sample(386)
        x =               26; #20833; // Sample(387)
        x =              236; #20833; // Sample(388)
        x =             -239; #20833; // Sample(389)
        x =               47; #20833; // Sample(390)
        x =             -262; #20833; // Sample(391)
        x =              214; #20833; // Sample(392)
        x =              156; #20833; // Sample(393)
        x =              229; #20833; // Sample(394)
        x =              102; #20833; // Sample(395)
        x =             -154; #20833; // Sample(396)
        x =              400; #20833; // Sample(397)
        x =              103; #20833; // Sample(398)
        x =              272; #20833; // Sample(399)
        x =              429; #20833; // Sample(400)
        x =              368; #20833; // Sample(401)
        x =              113; #20833; // Sample(402)
        x =              228; #20833; // Sample(403)
        x =              243; #20833; // Sample(404)
        x =              477; #20833; // Sample(405)
        x =              537; #20833; // Sample(406)
        x =               97; #20833; // Sample(407)
        x =              107; #20833; // Sample(408)
        x =              325; #20833; // Sample(409)
        x =              299; #20833; // Sample(410)
        x =              335; #20833; // Sample(411)
        x =               96; #20833; // Sample(412)
        x =               37; #20833; // Sample(413)
        x =              269; #20833; // Sample(414)
        x =              511; #20833; // Sample(415)
        x =              389; #20833; // Sample(416)
        x =              238; #20833; // Sample(417)
        x =              177; #20833; // Sample(418)
        x =               26; #20833; // Sample(419)
        x =              396; #20833; // Sample(420)
        x =              374; #20833; // Sample(421)
        x =              167; #20833; // Sample(422)
        x =              256; #20833; // Sample(423)
        x =              219; #20833; // Sample(424)
        x =              325; #20833; // Sample(425)
        x =              443; #20833; // Sample(426)
        x =             -217; #20833; // Sample(427)
        x =               38; #20833; // Sample(428)
        x =               63; #20833; // Sample(429)
        x =             -182; #20833; // Sample(430)
        x =              -16; #20833; // Sample(431)
        x =              174; #20833; // Sample(432)
        x =             -143; #20833; // Sample(433)
        x =             -417; #20833; // Sample(434)
        x =             -232; #20833; // Sample(435)
        x =               -5; #20833; // Sample(436)
        x =             -222; #20833; // Sample(437)
        x =               83; #20833; // Sample(438)
        x =             -220; #20833; // Sample(439)
        x =              -89; #20833; // Sample(440)
        x =             -263; #20833; // Sample(441)
        x =              -48; #20833; // Sample(442)
        x =             -493; #20833; // Sample(443)
        x =              112; #20833; // Sample(444)
        x =             -253; #20833; // Sample(445)
        x =             -252; #20833; // Sample(446)
        x =             -507; #20833; // Sample(447)
        x =             -249; #20833; // Sample(448)
        x =             -273; #20833; // Sample(449)
        x =             -497; #20833; // Sample(450)
        x =             -164; #20833; // Sample(451)
        x =               96; #20833; // Sample(452)
        x =              -65; #20833; // Sample(453)
        x =             -306; #20833; // Sample(454)
        x =             -192; #20833; // Sample(455)
        x =             -259; #20833; // Sample(456)
        x =             -221; #20833; // Sample(457)
        x =             -689; #20833; // Sample(458)
        x =             -468; #20833; // Sample(459)
        x =             -348; #20833; // Sample(460)
        x =             -170; #20833; // Sample(461)
        x =             -215; #20833; // Sample(462)
        x =             -296; #20833; // Sample(463)
        x =             -677; #20833; // Sample(464)
        x =             -529; #20833; // Sample(465)
        x =                4; #20833; // Sample(466)
        x =             -212; #20833; // Sample(467)
        x =             -223; #20833; // Sample(468)
        x =             -276; #20833; // Sample(469)
        x =              351; #20833; // Sample(470)
        x =             -312; #20833; // Sample(471)
        x =             -194; #20833; // Sample(472)
        x =              -49; #20833; // Sample(473)
        x =              117; #20833; // Sample(474)
        x =             -140; #20833; // Sample(475)
        x =               87; #20833; // Sample(476)
        x =              110; #20833; // Sample(477)
        x =              -10; #20833; // Sample(478)
        x =             -287; #20833; // Sample(479)
        x =              132; #20833; // Sample(480)
        x =               20; #20833; // Sample(481)
        x =              313; #20833; // Sample(482)
        x =             -119; #20833; // Sample(483)
        x =               58; #20833; // Sample(484)
        x =              -17; #20833; // Sample(485)
        x =             -251; #20833; // Sample(486)
        x =              -83; #20833; // Sample(487)
        x =             -236; #20833; // Sample(488)
        x =              469; #20833; // Sample(489)
        x =              213; #20833; // Sample(490)
        x =              296; #20833; // Sample(491)
        x =              237; #20833; // Sample(492)
        x =              423; #20833; // Sample(493)
        x =              512; #20833; // Sample(494)
        x =              162; #20833; // Sample(495)
        x =               67; #20833; // Sample(496)
        x =              469; #20833; // Sample(497)
        x =              693; #20833; // Sample(498)
        x =              236; #20833; // Sample(499)
        x =              141; #20833; // Sample(500)
        x =                0; #20833; // Sample(1)
        x =              183; #20833; // Sample(2)
        x =              290; #20833; // Sample(3)
        x =              277; #20833; // Sample(4)
        x =              150; #20833; // Sample(5)
        x =              -39; #20833; // Sample(6)
        x =             -212; #20833; // Sample(7)
        x =             -297; #20833; // Sample(8)
        x =             -260; #20833; // Sample(9)
        x =             -115; #20833; // Sample(10)
        x =               78; #20833; // Sample(11)
        x =              238; #20833; // Sample(12)
        x =              300; #20833; // Sample(13)
        x =              238; #20833; // Sample(14)
        x =               78; #20833; // Sample(15)
        x =             -115; #20833; // Sample(16)
        x =             -260; #20833; // Sample(17)
        x =             -297; #20833; // Sample(18)
        x =             -212; #20833; // Sample(19)
        x =              -39; #20833; // Sample(20)
        x =              150; #20833; // Sample(21)
        x =              277; #20833; // Sample(22)
        x =              290; #20833; // Sample(23)
        x =              183; #20833; // Sample(24)
        x =                0; #20833; // Sample(25)
        x =             -183; #20833; // Sample(26)
        x =             -290; #20833; // Sample(27)
        x =             -277; #20833; // Sample(28)
        x =             -150; #20833; // Sample(29)
        x =               39; #20833; // Sample(30)
        x =              212; #20833; // Sample(31)
        x =              297; #20833; // Sample(32)
        x =              260; #20833; // Sample(33)
        x =              115; #20833; // Sample(34)
        x =              -78; #20833; // Sample(35)
        x =             -238; #20833; // Sample(36)
        x =             -300; #20833; // Sample(37)
        x =             -238; #20833; // Sample(38)
        x =              -78; #20833; // Sample(39)
        x =              115; #20833; // Sample(40)
        x =              260; #20833; // Sample(41)
        x =              297; #20833; // Sample(42)
        x =              212; #20833; // Sample(43)
        x =               39; #20833; // Sample(44)
        x =             -150; #20833; // Sample(45)
        x =             -277; #20833; // Sample(46)
        x =             -290; #20833; // Sample(47)
        x =             -183; #20833; // Sample(48)
        x =               -0; #20833; // Sample(49)
        x =              183; #20833; // Sample(50)
        x =              290; #20833; // Sample(51)
        x =              277; #20833; // Sample(52)
        x =              150; #20833; // Sample(53)
        x =              -39; #20833; // Sample(54)
        x =             -212; #20833; // Sample(55)
        x =             -297; #20833; // Sample(56)
        x =             -260; #20833; // Sample(57)
        x =             -115; #20833; // Sample(58)
        x =               78; #20833; // Sample(59)
        x =              238; #20833; // Sample(60)
        x =              300; #20833; // Sample(61)
        x =              238; #20833; // Sample(62)
        x =               78; #20833; // Sample(63)
        x =             -115; #20833; // Sample(64)
        x =             -260; #20833; // Sample(65)
        x =             -297; #20833; // Sample(66)
        x =             -212; #20833; // Sample(67)
        x =              -39; #20833; // Sample(68)
        x =              150; #20833; // Sample(69)
        x =              277; #20833; // Sample(70)
        x =              290; #20833; // Sample(71)
        x =              183; #20833; // Sample(72)
        x =               -0; #20833; // Sample(73)
        x =             -183; #20833; // Sample(74)
        x =             -290; #20833; // Sample(75)
        x =             -277; #20833; // Sample(76)
        x =             -150; #20833; // Sample(77)
        x =               39; #20833; // Sample(78)
        x =              212; #20833; // Sample(79)
        x =              297; #20833; // Sample(80)
        x =              260; #20833; // Sample(81)
        x =              115; #20833; // Sample(82)
        x =              -78; #20833; // Sample(83)
        x =             -238; #20833; // Sample(84)
        x =             -300; #20833; // Sample(85)
        x =             -238; #20833; // Sample(86)
        x =              -78; #20833; // Sample(87)
        x =              115; #20833; // Sample(88)
        x =              260; #20833; // Sample(89)
        x =              297; #20833; // Sample(90)
        x =              212; #20833; // Sample(91)
        x =               39; #20833; // Sample(92)
        x =             -150; #20833; // Sample(93)
        x =             -277; #20833; // Sample(94)
        x =             -290; #20833; // Sample(95)
        x =             -183; #20833; // Sample(96)
        x =               -0; #20833; // Sample(97)
        x =              183; #20833; // Sample(98)
        x =              290; #20833; // Sample(99)
        x =              277; #20833; // Sample(100)
        x =              150; #20833; // Sample(101)
        x =              -39; #20833; // Sample(102)
        x =             -212; #20833; // Sample(103)
        x =             -297; #20833; // Sample(104)
        x =             -260; #20833; // Sample(105)
        x =             -115; #20833; // Sample(106)
        x =               78; #20833; // Sample(107)
        x =              238; #20833; // Sample(108)
        x =              300; #20833; // Sample(109)
        x =              238; #20833; // Sample(110)
        x =               78; #20833; // Sample(111)
        x =             -115; #20833; // Sample(112)
        x =             -260; #20833; // Sample(113)
        x =             -297; #20833; // Sample(114)
        x =             -212; #20833; // Sample(115)
        x =              -39; #20833; // Sample(116)
        x =              150; #20833; // Sample(117)
        x =              277; #20833; // Sample(118)
        x =              290; #20833; // Sample(119)
        x =              183; #20833; // Sample(120)
        x =               -0; #20833; // Sample(121)
        x =             -183; #20833; // Sample(122)
        x =             -290; #20833; // Sample(123)
        x =             -277; #20833; // Sample(124)
        x =             -150; #20833; // Sample(125)
        x =               39; #20833; // Sample(126)
        x =              212; #20833; // Sample(127)
        x =              297; #20833; // Sample(128)
        x =              260; #20833; // Sample(129)
        x =              115; #20833; // Sample(130)
        x =              -78; #20833; // Sample(131)
        x =             -238; #20833; // Sample(132)
        x =             -300; #20833; // Sample(133)
        x =             -238; #20833; // Sample(134)
        x =              -78; #20833; // Sample(135)
        x =              115; #20833; // Sample(136)
        x =              260; #20833; // Sample(137)
        x =              297; #20833; // Sample(138)
        x =              212; #20833; // Sample(139)
        x =               39; #20833; // Sample(140)
        x =             -150; #20833; // Sample(141)
        x =             -277; #20833; // Sample(142)
        x =             -290; #20833; // Sample(143)
        x =             -183; #20833; // Sample(144)
        x =                0; #20833; // Sample(145)
        x =              183; #20833; // Sample(146)
        x =              290; #20833; // Sample(147)
        x =              277; #20833; // Sample(148)
        x =              150; #20833; // Sample(149)
        x =              -39; #20833; // Sample(150)
        x =             -212; #20833; // Sample(151)
        x =             -297; #20833; // Sample(152)
        x =             -260; #20833; // Sample(153)
        x =             -115; #20833; // Sample(154)
        x =               78; #20833; // Sample(155)
        x =              238; #20833; // Sample(156)
        x =              300; #20833; // Sample(157)
        x =              238; #20833; // Sample(158)
        x =               78; #20833; // Sample(159)
        x =             -115; #20833; // Sample(160)
        x =             -260; #20833; // Sample(161)
        x =             -297; #20833; // Sample(162)
        x =             -212; #20833; // Sample(163)
        x =              -39; #20833; // Sample(164)
        x =              150; #20833; // Sample(165)
        x =              277; #20833; // Sample(166)
        x =              290; #20833; // Sample(167)
        x =              183; #20833; // Sample(168)
        x =               -0; #20833; // Sample(169)
        x =             -183; #20833; // Sample(170)
        x =             -290; #20833; // Sample(171)
        x =             -277; #20833; // Sample(172)
        x =             -150; #20833; // Sample(173)
        x =               39; #20833; // Sample(174)
        x =              212; #20833; // Sample(175)
        x =              297; #20833; // Sample(176)
        x =              260; #20833; // Sample(177)
        x =              115; #20833; // Sample(178)
        x =              -78; #20833; // Sample(179)
        x =             -238; #20833; // Sample(180)
        x =             -300; #20833; // Sample(181)
        x =             -238; #20833; // Sample(182)
        x =              -78; #20833; // Sample(183)
        x =              115; #20833; // Sample(184)
        x =              260; #20833; // Sample(185)
        x =              297; #20833; // Sample(186)
        x =              212; #20833; // Sample(187)
        x =               39; #20833; // Sample(188)
        x =             -150; #20833; // Sample(189)
        x =             -277; #20833; // Sample(190)
        x =             -290; #20833; // Sample(191)
        x =             -183; #20833; // Sample(192)
        x =               -0; #20833; // Sample(193)
        x =              183; #20833; // Sample(194)
        x =              290; #20833; // Sample(195)
        x =              277; #20833; // Sample(196)
        x =              150; #20833; // Sample(197)
        x =              -39; #20833; // Sample(198)
        x =             -212; #20833; // Sample(199)
        x =             -297; #20833; // Sample(200)
        x =             -260; #20833; // Sample(201)
        x =             -115; #20833; // Sample(202)
        x =               78; #20833; // Sample(203)
        x =              238; #20833; // Sample(204)
        x =              300; #20833; // Sample(205)
        x =              238; #20833; // Sample(206)
        x =               78; #20833; // Sample(207)
        x =             -115; #20833; // Sample(208)
        x =             -260; #20833; // Sample(209)
        x =             -297; #20833; // Sample(210)
        x =             -212; #20833; // Sample(211)
        x =              -39; #20833; // Sample(212)
        x =              150; #20833; // Sample(213)
        x =              277; #20833; // Sample(214)
        x =              290; #20833; // Sample(215)
        x =              183; #20833; // Sample(216)
        x =                0; #20833; // Sample(217)
        x =             -183; #20833; // Sample(218)
        x =             -290; #20833; // Sample(219)
        x =             -277; #20833; // Sample(220)
        x =             -150; #20833; // Sample(221)
        x =               39; #20833; // Sample(222)
        x =              212; #20833; // Sample(223)
        x =              297; #20833; // Sample(224)
        x =              260; #20833; // Sample(225)
        x =              115; #20833; // Sample(226)
        x =              -78; #20833; // Sample(227)
        x =             -238; #20833; // Sample(228)
        x =             -300; #20833; // Sample(229)
        x =             -238; #20833; // Sample(230)
        x =              -78; #20833; // Sample(231)
        x =              115; #20833; // Sample(232)
        x =              260; #20833; // Sample(233)
        x =              297; #20833; // Sample(234)
        x =              212; #20833; // Sample(235)
        x =               39; #20833; // Sample(236)
        x =             -150; #20833; // Sample(237)
        x =             -277; #20833; // Sample(238)
        x =             -290; #20833; // Sample(239)
        x =             -183; #20833; // Sample(240)
        x =                0; #20833; // Sample(241)
        x =              183; #20833; // Sample(242)
        x =              290; #20833; // Sample(243)
        x =              277; #20833; // Sample(244)
        x =              150; #20833; // Sample(245)
        x =              -39; #20833; // Sample(246)
        x =             -212; #20833; // Sample(247)
        x =             -297; #20833; // Sample(248)
        x =             -260; #20833; // Sample(249)
        x =             -115; #20833; // Sample(250)
        x =               78; #20833; // Sample(251)
        x =              238; #20833; // Sample(252)
        x =              300; #20833; // Sample(253)
        x =              238; #20833; // Sample(254)
        x =               78; #20833; // Sample(255)
        x =             -115; #20833; // Sample(256)
        x =             -260; #20833; // Sample(257)
        x =             -297; #20833; // Sample(258)
        x =             -212; #20833; // Sample(259)
        x =              -39; #20833; // Sample(260)
        x =              150; #20833; // Sample(261)
        x =              277; #20833; // Sample(262)
        x =              290; #20833; // Sample(263)
        x =              183; #20833; // Sample(264)
        x =               -0; #20833; // Sample(265)
        x =             -183; #20833; // Sample(266)
        x =             -290; #20833; // Sample(267)
        x =             -277; #20833; // Sample(268)
        x =             -150; #20833; // Sample(269)
        x =               39; #20833; // Sample(270)
        x =              212; #20833; // Sample(271)
        x =              297; #20833; // Sample(272)
        x =              260; #20833; // Sample(273)
        x =              115; #20833; // Sample(274)
        x =              -78; #20833; // Sample(275)
        x =             -238; #20833; // Sample(276)
        x =             -300; #20833; // Sample(277)
        x =             -238; #20833; // Sample(278)
        x =              -78; #20833; // Sample(279)
        x =              115; #20833; // Sample(280)
        x =              260; #20833; // Sample(281)
        x =              297; #20833; // Sample(282)
        x =              212; #20833; // Sample(283)
        x =               39; #20833; // Sample(284)
        x =             -150; #20833; // Sample(285)
        x =             -277; #20833; // Sample(286)
        x =             -290; #20833; // Sample(287)
        x =             -183; #20833; // Sample(288)
        x =                0; #20833; // Sample(289)
        x =              183; #20833; // Sample(290)
        x =              290; #20833; // Sample(291)
        x =              277; #20833; // Sample(292)
        x =              150; #20833; // Sample(293)
        x =              -39; #20833; // Sample(294)
        x =             -212; #20833; // Sample(295)
        x =             -297; #20833; // Sample(296)
        x =             -260; #20833; // Sample(297)
        x =             -115; #20833; // Sample(298)
        x =               78; #20833; // Sample(299)
        x =              238; #20833; // Sample(300)
        x =              300; #20833; // Sample(301)
        x =              238; #20833; // Sample(302)
        x =               78; #20833; // Sample(303)
        x =             -115; #20833; // Sample(304)
        x =             -260; #20833; // Sample(305)
        x =             -297; #20833; // Sample(306)
        x =             -212; #20833; // Sample(307)
        x =              -39; #20833; // Sample(308)
        x =              150; #20833; // Sample(309)
        x =              277; #20833; // Sample(310)
        x =              290; #20833; // Sample(311)
        x =              183; #20833; // Sample(312)
        x =               -0; #20833; // Sample(313)
        x =             -183; #20833; // Sample(314)
        x =             -290; #20833; // Sample(315)
        x =             -277; #20833; // Sample(316)
        x =             -150; #20833; // Sample(317)
        x =               39; #20833; // Sample(318)
        x =              212; #20833; // Sample(319)
        x =              297; #20833; // Sample(320)
        x =              260; #20833; // Sample(321)
        x =              115; #20833; // Sample(322)
        x =              -78; #20833; // Sample(323)
        x =             -238; #20833; // Sample(324)
        x =             -300; #20833; // Sample(325)
        x =             -238; #20833; // Sample(326)
        x =              -78; #20833; // Sample(327)
        x =              115; #20833; // Sample(328)
        x =              260; #20833; // Sample(329)
        x =              297; #20833; // Sample(330)
        x =              212; #20833; // Sample(331)
        x =               39; #20833; // Sample(332)
        x =             -150; #20833; // Sample(333)
        x =             -277; #20833; // Sample(334)
        x =             -290; #20833; // Sample(335)
        x =             -183; #20833; // Sample(336)
        x =                0; #20833; // Sample(337)
        x =              183; #20833; // Sample(338)
        x =              290; #20833; // Sample(339)
        x =              277; #20833; // Sample(340)
        x =              150; #20833; // Sample(341)
        x =              -39; #20833; // Sample(342)
        x =             -212; #20833; // Sample(343)
        x =             -297; #20833; // Sample(344)
        x =             -260; #20833; // Sample(345)
        x =             -115; #20833; // Sample(346)
        x =               78; #20833; // Sample(347)
        x =              238; #20833; // Sample(348)
        x =              300; #20833; // Sample(349)
        x =              238; #20833; // Sample(350)
        x =               78; #20833; // Sample(351)
        x =             -115; #20833; // Sample(352)
        x =             -260; #20833; // Sample(353)
        x =             -297; #20833; // Sample(354)
        x =             -212; #20833; // Sample(355)
        x =              -39; #20833; // Sample(356)
        x =              150; #20833; // Sample(357)
        x =              277; #20833; // Sample(358)
        x =              290; #20833; // Sample(359)
        x =              183; #20833; // Sample(360)
        x =               -0; #20833; // Sample(361)
        x =             -183; #20833; // Sample(362)
        x =             -290; #20833; // Sample(363)
        x =             -277; #20833; // Sample(364)
        x =             -150; #20833; // Sample(365)
        x =               39; #20833; // Sample(366)
        x =              212; #20833; // Sample(367)
        x =              297; #20833; // Sample(368)
        x =              260; #20833; // Sample(369)
        x =              115; #20833; // Sample(370)
        x =              -78; #20833; // Sample(371)
        x =             -238; #20833; // Sample(372)
        x =             -300; #20833; // Sample(373)
        x =             -238; #20833; // Sample(374)
        x =              -78; #20833; // Sample(375)
        x =              115; #20833; // Sample(376)
        x =              260; #20833; // Sample(377)
        x =              297; #20833; // Sample(378)
        x =              212; #20833; // Sample(379)
        x =               39; #20833; // Sample(380)
        x =             -150; #20833; // Sample(381)
        x =             -277; #20833; // Sample(382)
        x =             -290; #20833; // Sample(383)
        x =             -183; #20833; // Sample(384)
        x =               -0; #20833; // Sample(385)
        x =              183; #20833; // Sample(386)
        x =              290; #20833; // Sample(387)
        x =              277; #20833; // Sample(388)
        x =              150; #20833; // Sample(389)
        x =              -39; #20833; // Sample(390)
        x =             -212; #20833; // Sample(391)
        x =             -297; #20833; // Sample(392)
        x =             -260; #20833; // Sample(393)
        x =             -115; #20833; // Sample(394)
        x =               78; #20833; // Sample(395)
        x =              238; #20833; // Sample(396)
        x =              300; #20833; // Sample(397)
        x =              238; #20833; // Sample(398)
        x =               78; #20833; // Sample(399)
        x =             -115; #20833; // Sample(400)
        x =             -260; #20833; // Sample(401)
        x =             -297; #20833; // Sample(402)
        x =             -212; #20833; // Sample(403)
        x =              -39; #20833; // Sample(404)
        x =              150; #20833; // Sample(405)
        x =              277; #20833; // Sample(406)
        x =              290; #20833; // Sample(407)
        x =              183; #20833; // Sample(408)
        x =                0; #20833; // Sample(409)
        x =             -183; #20833; // Sample(410)
        x =             -290; #20833; // Sample(411)
        x =             -277; #20833; // Sample(412)
        x =             -150; #20833; // Sample(413)
        x =               39; #20833; // Sample(414)
        x =              212; #20833; // Sample(415)
        x =              297; #20833; // Sample(416)
        x =              260; #20833; // Sample(417)
        x =              115; #20833; // Sample(418)
        x =              -78; #20833; // Sample(419)
        x =             -238; #20833; // Sample(420)
        x =             -300; #20833; // Sample(421)
        x =             -238; #20833; // Sample(422)
        x =              -78; #20833; // Sample(423)
        x =              115; #20833; // Sample(424)
        x =              260; #20833; // Sample(425)
        x =              297; #20833; // Sample(426)
        x =              212; #20833; // Sample(427)
        x =               39; #20833; // Sample(428)
        x =             -150; #20833; // Sample(429)
        x =             -277; #20833; // Sample(430)
        x =             -290; #20833; // Sample(431)
        x =             -183; #20833; // Sample(432)
        x =               -0; #20833; // Sample(433)
        x =              183; #20833; // Sample(434)
        x =              290; #20833; // Sample(435)
        x =              277; #20833; // Sample(436)
        x =              150; #20833; // Sample(437)
        x =              -39; #20833; // Sample(438)
        x =             -212; #20833; // Sample(439)
        x =             -297; #20833; // Sample(440)
        x =             -260; #20833; // Sample(441)
        x =             -115; #20833; // Sample(442)
        x =               78; #20833; // Sample(443)
        x =              238; #20833; // Sample(444)
        x =              300; #20833; // Sample(445)
        x =              238; #20833; // Sample(446)
        x =               78; #20833; // Sample(447)
        x =             -115; #20833; // Sample(448)
        x =             -260; #20833; // Sample(449)
        x =             -297; #20833; // Sample(450)
        x =             -212; #20833; // Sample(451)
        x =              -39; #20833; // Sample(452)
        x =              150; #20833; // Sample(453)
        x =              277; #20833; // Sample(454)
        x =              290; #20833; // Sample(455)
        x =              183; #20833; // Sample(456)
        x =                0; #20833; // Sample(457)
        x =             -183; #20833; // Sample(458)
        x =             -290; #20833; // Sample(459)
        x =             -277; #20833; // Sample(460)
        x =             -150; #20833; // Sample(461)
        x =               39; #20833; // Sample(462)
        x =              212; #20833; // Sample(463)
        x =              297; #20833; // Sample(464)
        x =              260; #20833; // Sample(465)
        x =              115; #20833; // Sample(466)
        x =              -78; #20833; // Sample(467)
        x =             -238; #20833; // Sample(468)
        x =             -300; #20833; // Sample(469)
        x =             -238; #20833; // Sample(470)
        x =              -78; #20833; // Sample(471)
        x =              115; #20833; // Sample(472)
        x =              260; #20833; // Sample(473)
        x =              297; #20833; // Sample(474)
        x =              212; #20833; // Sample(475)
        x =               39; #20833; // Sample(476)
        x =             -150; #20833; // Sample(477)
        x =             -277; #20833; // Sample(478)
        x =             -290; #20833; // Sample(479)
        x =             -183; #20833; // Sample(480)
        x =                0; #20833; // Sample(481)
        x =              183; #20833; // Sample(482)
        x =              290; #20833; // Sample(483)
        x =              277; #20833; // Sample(484)
        x =              150; #20833; // Sample(485)
        x =              -39; #20833; // Sample(486)
        x =             -212; #20833; // Sample(487)
        x =             -297; #20833; // Sample(488)
        x =             -260; #20833; // Sample(489)
        x =             -115; #20833; // Sample(490)
        x =               78; #20833; // Sample(491)
        x =              238; #20833; // Sample(492)
        x =              300; #20833; // Sample(493)
        x =              238; #20833; // Sample(494)
        x =               78; #20833; // Sample(495)
        x =             -115; #20833; // Sample(496)
        x =             -260; #20833; // Sample(497)
        x =             -297; #20833; // Sample(498)
        x =             -212; #20833; // Sample(499)
        x =              -39; #20833; // Sample(500)
        $stop;
    end
endmodule
